///////////////////////////////////////////////////////////////////////////////
// File: usb_hid_keyboard_engine.v (FIXED VERSION)
// Description: USB HID Keyboard Host Engine
//
// FIXES APPLIED:
// - CRITICAL: Added missing 'end' statement to close STATE_WAIT_SOF
// - CRITICAL: Fixed array indexing - rx_buffer is packed, not unpacked
// - CRITICAL: Changed rx_count from [3:0] to [6:0] to support 64 bytes
// - Simplified report packing (removed 64-iteration for loop)
// - Now uses wire definitions for byte extraction
//
// Polls a USB HID keyboard device for keypress data via interrupt endpoint.
// Supports both Boot Protocol (8 bytes) and Report Protocol (variable length).
///////////////////////////////////////////////////////////////////////////////

module usb_hid_keyboard_engine (
    // Clock and Reset
    input  wire        clk,
    input  wire        rst_n,
    
    // Control Interface
    input  wire        enable,
    input  wire        enumerated,
    
    // Device Information
    input  wire [6:0]  device_addr,
    input  wire [3:0]  endp_number,
    input  wire [7:0]  max_packet_size,
    input  wire [1:0]  device_speed,
    input  wire [7:0]  poll_interval,
    
    // Token Generator Interface
    output reg         token_start,
    output reg  [1:0]  token_type,
    output reg  [6:0]  token_addr,
    output reg  [3:0]  token_endp,
    input  wire        token_ready,
    input  wire        token_done,
    
    // UTMI Receive Interface
    input  wire [7:0]  utmi_rx_data,
    input  wire        utmi_rx_valid,
    input  wire        utmi_rx_active,
    input  wire [3:0]  utmi_rx_pid,
    
    // SOF Interface
    input  wire        sof_trigger,
    input  wire [10:0] frame_number,
    
    // Keyboard Report Output
    output reg         report_valid,
    output reg  [63:0] report_data,
    output reg  [6:0]  report_length,
    
    // Decoded Boot Protocol Fields
    output reg  [7:0]  report_modifiers,
    output reg  [7:0]  report_key0,
    output reg  [7:0]  report_key1,
    output reg  [7:0]  report_key2,
    output reg  [7:0]  report_key3,
    output reg  [7:0]  report_key4,
    output reg  [7:0]  report_key5,
    
    // Status
    output reg  [7:0]  status,
    output reg  [15:0] poll_count,
    output reg         active           // Polling activity indicator
);

    // Token types
    localparam TOKEN_IN = 2'b01;
    
    // Speed definitions
    localparam SPEED_LOW = 2'b00;
    localparam SPEED_FULL = 2'b01;
    localparam SPEED_HIGH = 2'b10;
    
    // PIDs
    localparam PID_DATA0 = 4'b0011;
    localparam PID_DATA1 = 4'b1011;
    localparam PID_ACK   = 4'b0010;
    localparam PID_NAK   = 4'b1010;
    localparam PID_STALL = 4'b1110;
    
    // State Machine
    localparam STATE_IDLE           = 3'd0;
    localparam STATE_WAIT_SOF       = 3'd1;
    localparam STATE_SEND_IN_TOKEN  = 3'd2;
    localparam STATE_WAIT_DATA      = 3'd3;
    localparam STATE_PROCESS_DATA   = 3'd4;
    localparam STATE_SEND_ACK       = 3'd5;
    localparam STATE_ERROR          = 3'd6;
    
    reg [2:0]  state;
    reg [63:0] rx_buffer;
    reg [6:0]  rx_count;            // FIXED: Changed from [3:0] to [6:0]
    reg        data_pid;
    
    // Byte accessors for packed buffer
    wire [7:0] rx_byte0 = rx_buffer[7:0];
    wire [7:0] rx_byte1 = rx_buffer[15:8];
    wire [7:0] rx_byte2 = rx_buffer[23:16];
    wire [7:0] rx_byte3 = rx_buffer[31:24];
    wire [7:0] rx_byte4 = rx_buffer[39:32];
    wire [7:0] rx_byte5 = rx_buffer[47:40];
    wire [7:0] rx_byte6 = rx_buffer[55:48];
    wire [7:0] rx_byte7 = rx_buffer[63:56];
    
    reg [10:0] last_frame;
    reg [7:0]  poll_counter;
    reg [7:0]  effective_interval;
    reg [31:0] timeout_counter;
    reg [3:0]  error_count;
    reg [31:0] watchdog_counter;
    
    // Watchdog timeout: 3 seconds at 60MHz
    localparam WATCHDOG_TIMEOUT = 32'd180000000;
    
    // Status bits
    localparam STATUS_ACTIVE     = 8'h01;
    localparam STATUS_ERROR      = 8'h02;
    localparam STATUS_STALL      = 8'h04;
    localparam STATUS_TIMEOUT    = 8'h08;
    localparam STATUS_ENUMERATED = 8'h10;
    
    integer i;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= STATE_IDLE;
            token_start <= 1'b0;
            token_type <= 2'd0;
            token_addr <= 7'd0;
            token_endp <= 4'd0;
            report_valid <= 1'b0;
            report_data <= 512'd0;
            report_length <= 7'd0;
            report_modifiers <= 8'd0;
            report_key0 <= 8'd0;
            report_key1 <= 8'd0;
            report_key2 <= 8'd0;
            report_key3 <= 8'd0;
            report_key4 <= 8'd0;
            report_key5 <= 8'd0;
            status <= 8'd0;
            poll_count <= 16'd0;
            active <= 1'b0;
            rx_count <= 7'd0;
            data_pid <= 1'b0;
            last_frame <= 11'd0;
            poll_counter <= 8'd0;
            effective_interval <= 8'd1;
            timeout_counter <= 32'd0;
            error_count <= 4'd0;
            watchdog_counter <= 32'd0;
            rx_buffer <= 64'd0;
        end else begin
            // Default outputs
            token_start <= 1'b0;
            report_valid <= 1'b0;
            active <= (state != STATE_IDLE) && enable && enumerated;
            
            // Watchdog counter
            if (state != STATE_IDLE && enable && enumerated)
                watchdog_counter <= watchdog_counter + 1'b1;
            else
                watchdog_counter <= 32'd0;
            
            // Watchdog timeout
            if (watchdog_counter >= WATCHDOG_TIMEOUT) begin
                state <= STATE_IDLE;
                status <= STATUS_TIMEOUT;
                watchdog_counter <= 32'd0;
            end
            
            // FIXED: Collect RX data using shift register
            if (utmi_rx_valid && rx_count < 7'd8) begin
                rx_buffer <= {utmi_rx_data, rx_buffer[63:8]};
                rx_count <= rx_count + 1'b1;
            end
            
            // Timeout counter
            timeout_counter <= timeout_counter + 1'b1;
            
            case (state)
                STATE_IDLE: begin
                    status <= enumerated ? STATUS_ENUMERATED : 8'h00;
                    timeout_counter <= 32'd0;
                    error_count <= 4'd0;
                    
                    if (enable && enumerated) begin
                        state <= STATE_WAIT_SOF;
                        data_pid <= 1'b0;
                    end
                end
                
                STATE_WAIT_SOF: begin
                    status <= STATUS_ACTIVE | STATUS_ENUMERATED;
                    
                    if (sof_trigger && frame_number != last_frame) begin
                        last_frame <= frame_number;
                        
                        // Calculate effective interval based on speed
                        if (device_speed == SPEED_HIGH) begin
                            // Limit shift to prevent overflow
                            if (poll_interval > 8'd8)
                                effective_interval <= 8'd128;
                            else
                                effective_interval <= (8'd1 << (poll_interval - 1));
                        end else begin
                            effective_interval <= poll_interval;
                        end
                        
                        if (poll_counter >= effective_interval - 1) begin
                            poll_counter <= 8'd0;
                            rx_count <= 7'd0;
                            state <= STATE_SEND_IN_TOKEN;
                            timeout_counter <= 32'd0;
                            watchdog_counter <= 32'd0;
                        end else begin
                            poll_counter <= poll_counter + 1'b1;
                        end
                    end
                end  // FIXED: Added missing 'end' to close STATE_WAIT_SOF
                
                STATE_SEND_IN_TOKEN: begin
                    if (token_ready && !token_start) begin
                        token_start <= 1'b1;
                        token_type <= TOKEN_IN;
                        token_addr <= device_addr;
                        token_endp <= endp_number;
                        state <= STATE_WAIT_DATA;
                        timeout_counter <= 32'd0;
                    end
                end
                
                STATE_WAIT_DATA: begin
                    if (!utmi_rx_active && rx_count > 7'd0) begin
                        if ((data_pid == 1'b0 && utmi_rx_pid == PID_DATA0) ||
                            (data_pid == 1'b1 && utmi_rx_pid == PID_DATA1)) begin
                            state <= STATE_PROCESS_DATA;
                            watchdog_counter <= 32'd0;
                        end else if (utmi_rx_pid == PID_NAK) begin
                            state <= STATE_WAIT_SOF;
                            watchdog_counter <= 32'd0;
                        end else if (utmi_rx_pid == PID_STALL) begin
                            status <= STATUS_STALL;
                            error_count <= error_count + 1'b1;
                            state <= STATE_ERROR;
                        end
                    end
                    
                    // Timeout after 10ms
                    if (timeout_counter > 32'd600000) begin
                        error_count <= error_count + 1'b1;
                        if (error_count >= 4'd10) begin
                            status <= STATUS_TIMEOUT;
                            state <= STATE_ERROR;
                        end else begin
                            state <= STATE_WAIT_SOF;
                        end
                    end
                end
                
                STATE_PROCESS_DATA: begin
                    if (rx_count >= 7'd3) begin
                        // FIXED: Simplified report packing using wire definitions
                        report_data[7:0]    <= rx_byte0;
                        report_data[15:8]   <= (rx_count > 7'd1) ? rx_byte1 : 8'd0;
                        report_data[23:16]  <= (rx_count > 7'd2) ? rx_byte2 : 8'd0;
                        report_data[31:24]  <= (rx_count > 7'd3) ? rx_byte3 : 8'd0;
                        report_data[39:32]  <= (rx_count > 7'd4) ? rx_byte4 : 8'd0;
                        report_data[47:40]  <= (rx_count > 7'd5) ? rx_byte5 : 8'd0;
                        report_data[55:48]  <= (rx_count > 7'd6) ? rx_byte6 : 8'd0;
                        report_data[63:56]  <= (rx_count > 7'd7) ? rx_byte7 : 8'd0;
                        // Note: report_data is only 64 bits, removed invalid [511:64] assignment
                        
                        report_length <= rx_count;
                        
                        // FIXED: Decode boot protocol using wire definitions
                        if (rx_count >= 7'd8) begin
                            report_modifiers <= rx_byte0;
                            // rx_byte1 is reserved in boot protocol
                            report_key0 <= rx_byte2;
                            report_key1 <= rx_byte3;
                            report_key2 <= rx_byte4;
                            report_key3 <= rx_byte5;
                            report_key4 <= rx_byte6;
                            report_key5 <= rx_byte7;
                        end else begin
                            report_modifiers <= rx_byte0;
                            report_key0 <= (rx_count > 7'd1) ? rx_byte1 : 8'd0;
                            report_key1 <= (rx_count > 7'd2) ? rx_byte2 : 8'd0;
                            report_key2 <= (rx_count > 7'd3) ? rx_byte3 : 8'd0;
                            report_key3 <= (rx_count > 7'd4) ? rx_byte4 : 8'd0;
                            report_key4 <= (rx_count > 7'd5) ? rx_byte5 : 8'd0;
                            report_key5 <= (rx_count > 7'd6) ? rx_byte6 : 8'd0;
                        end
                        
                        report_valid <= 1'b1;
                        data_pid <= ~data_pid;
                        poll_count <= poll_count + 1'b1;
                    end
                    
                    state <= STATE_WAIT_SOF;
                end
                
                STATE_ERROR: begin
                    if (!enable) begin
                        state <= STATE_IDLE;
                    end
                end
                
                default: state <= STATE_IDLE;
            endcase
        end
    end

endmodule