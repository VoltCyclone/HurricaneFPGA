///////////////////////////////////////////////////////////////////////////////
// File: usb_phy_wrapper.v (FIXED VERSION)
// Description: USB PHY interface wrapper for ECP5 FPGA
//
// FIXES APPLIED:
// - CRITICAL: Added proper CDC synchronizer chain for line_state crossing
//   from clk domain to clk_480mhz domain (2-flop synchronizer)
// - CRITICAL: Removed combinatorial clock (clk_recovered) - now using it as
//   clock enable with edge detection instead
// - Fixed metastability risk in bit_phase_detector
// - Fixed EOP detection to use synchronized line state
//
// This module provides a wrapper for the USB physical interfaces, handling the
// low-level signaling for USB 2.0 data transmission and reception.
//
// Target: Lattice ECP5 on Cynthion device
///////////////////////////////////////////////////////////////////////////////

module usb_phy_wrapper (
    // Clock and Reset
    input  wire       clk,              // System clock (60MHz)
    input  wire       clk_480mhz,       // High-speed bit clock (480MHz)
    input  wire       rst_n,            // Active low reset

    // PHY Interface Pins
    input  wire       usb_dp_i,         // USB D+ input
    input  wire       usb_dn_i,         // USB D- input
    output wire       usb_dp_o,         // USB D+ output
    output wire       usb_dn_o,         // USB D- output
    output wire       usb_dp_oe,        // USB D+ output enable
    output wire       usb_dn_oe,        // USB D- output enable
    output wire       usb_pullup_en,    // USB pull-up resistor enable

    // UTMI Interface
    output wire [1:0] utmi_line_state,  // USB line state (SE0, J, K, SE1)
    output wire [7:0] utmi_rx_data,     // Received data
    output wire       utmi_rx_valid,    // Received data valid
    output wire       utmi_rx_active,   // Receiving packet
    output wire       utmi_rx_error,    // Receive error
    input  wire [7:0] utmi_tx_data,     // Data to transmit
    input  wire       utmi_tx_valid,    // Data valid for transmission
    output wire       utmi_tx_ready,    // PHY ready for transmission
    input  wire [1:0] utmi_tx_op_mode,  // Transmit operation mode
    input  wire [1:0] utmi_xcvr_select, // Transceiver speed selection
    input  wire       utmi_termselect,  // Termination selection
    input  wire       utmi_dppulldown,  // D+ pulldown enable
    input  wire       utmi_dmpulldown,  // D- pulldown enable
    
    // PHY Monitoring Interface (for debug)
    output wire [1:0] phy_line_state,   // Current raw line state for monitoring
    output wire       phy_rx_carrier,   // Carrier detect
    output wire       phy_rx_clock,     // Recovered clock
    
    // Configuration and Control
    input  wire [1:0] usb_speed_ctrl,   // USB speed selection (00=LS, 01=FS, 10=HS)
    input  wire       phy_reset,        // PHY-specific reset
    output wire       phy_status        // PHY status (connected, speed, etc.)
);

    // Internal signals
    reg  [1:0]  line_state_q;           // Registered line state (clk domain)
    reg  [1:0]  line_state_sync;        // Synchronized line state
    
    // ADDED: CDC synchronizer chain for clk_480mhz domain
    reg  [1:0]  line_state_480_sync1;   // First stage synchronizer
    reg  [1:0]  line_state_480_sync2;   // Second stage synchronizer
    
    reg  [7:0]  shift_reg;              // NRZI bit shift register
    reg         bit_phase_detector;     // Phase detection for clock recovery
    reg         bit_stuff_counter;      // Bit stuffing counter
    reg         rx_active_r;            // Registered rx_active
    reg         tx_busy;                // Transmitter busy flag
    
    // ADDED: Clock enable edge detection
    reg         clk_recovered_prev;
    wire        clk_recovered_edge;
    
    wire        nrzi_data;              // NRZI encoded outgoing data
    wire        clk_recovered;          // Clock recovery signal (used as enable, not clock)
    wire        sync_detect;            // SYNC pattern detection
    wire        eop_detect;             // End of packet detection

    // NRZI encoding/decoding logic
    // ----------------------------

    // Line state synchronization
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            line_state_q <= 2'b00;
            line_state_sync <= 2'b00;
        end else begin
            line_state_sync <= {usb_dn_i, usb_dp_i};
            line_state_q <= line_state_sync;
        end
    end

    // Assign the UTMI line state
    assign utmi_line_state = line_state_q;
    
    // Assign the raw line state for monitoring
    assign phy_line_state = line_state_q;

    // Clock recovery and NRZI decoding
    // -------------------------------
    // FIXED: Added proper CDC and removed combinatorial clock
    // For accurate implementation, we need complex CDR (Clock Data Recovery)
    // The simplified version below would be expanded in a real implementation

    // FIXED: CDC synchronizer chain from clk to clk_480mhz domain
    always @(posedge clk_480mhz or negedge rst_n) begin
        if (!rst_n) begin
            line_state_480_sync1 <= 2'b00;
            line_state_480_sync2 <= 2'b00;
        end else begin
            line_state_480_sync1 <= line_state_q;         // First flop
            line_state_480_sync2 <= line_state_480_sync1; // Second flop - safe to use
        end
    end

    // Detect transitions for clock recovery using SYNCHRONIZED line state
    always @(posedge clk_480mhz or negedge rst_n) begin
        if (!rst_n) begin
            bit_phase_detector <= 1'b0;
            rx_active_r <= 1'b0;
        end else begin
            bit_phase_detector <= line_state_480_sync2[0] ^ line_state_480_sync2[1]; // Use synchronized version
            rx_active_r <= sync_detect | (rx_active_r & ~eop_detect);
        end
    end

    // Simplified CDR implementation (used as enable, not clock)
    assign clk_recovered = bit_phase_detector & rx_active_r;
    assign clk_recovered_edge = clk_recovered & ~clk_recovered_prev;
    assign phy_rx_clock = clk_recovered; // For monitoring
    
    // SYNC pattern detection (simplified)
    assign sync_detect = (shift_reg == 8'b10000000); // SYNC = K J K J K J K K
    
    // EOP detection (simplified) - use synchronized line state
    assign eop_detect = (line_state_480_sync2 == 2'b00) & rx_active_r; // SE0 condition
    
    // FIXED: Use proper clock with enable instead of combinatorial clock
    always @(posedge clk_480mhz or negedge rst_n) begin
        if (!rst_n) begin
            shift_reg <= 8'h00;
            clk_recovered_prev <= 1'b0;
        end else begin
            clk_recovered_prev <= clk_recovered;
            
            // Only shift on rising edge of recovered clock
            if (clk_recovered_edge && rx_active_r) begin
                // NRZI decoding and bit stuffing removal would be implemented here
                shift_reg <= {shift_reg[6:0], line_state_480_sync2[0]};
            end
        end
    end

    // Transmitter logic
    // ----------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            tx_busy <= 1'b0;
        end else begin
            if (utmi_tx_valid && !tx_busy) begin
                tx_busy <= 1'b1;
            end else if (!utmi_tx_valid) begin
                tx_busy <= 1'b0;
            end
        end
    end
    
    // NRZI encoding for transmission (simplified)
    // In real implementation, would include bit stuffing and full NRZI processing
    assign nrzi_data = utmi_tx_valid ? utmi_tx_data[0] : 1'b1; // Idle = J state
    
    // Output assignments
    assign usb_dp_o = (utmi_tx_op_mode == 2'b00) ? 1'b1 : nrzi_data;
    assign usb_dn_o = (utmi_tx_op_mode == 2'b00) ? 1'b0 : ~nrzi_data;
    assign usb_dp_oe = tx_busy;
    assign usb_dn_oe = tx_busy;
    
    // Pull-up resistor control based on speed and mode
    assign usb_pullup_en = (utmi_xcvr_select != 2'b00);
    
    // Assign UTMI Rx signals (simplified - full implementation would need proper DPLL)
    assign utmi_rx_data = shift_reg;
    assign utmi_rx_valid = rx_active_r & ~(|shift_reg[1:0]); // Simplified data valid check
    assign utmi_rx_active = rx_active_r;
    assign utmi_rx_error = rx_active_r & eop_detect & (shift_reg[7:0] != 8'h00); // Simplified error detection
    
    // Transmit ready signal
    assign utmi_tx_ready = ~tx_busy;
    
    // Carrier detection (simplified)
    assign phy_rx_carrier = (utmi_line_state != 2'b00);
    
    // PHY status - in a real implementation, this would report negotiated speed, connection status, etc.
    assign phy_status = (utmi_line_state != 2'b00); // Simplified - just check if non-SE0

endmodule